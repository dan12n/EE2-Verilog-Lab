module add3_ge5 (in, out); //W1 is input, and A1 is output
	input [3:0] in;
	output [3:0] out;

	reg [3:0] out;
	
	always @(*)
		case (in)
		//IF not greater than five
		 4'b0000: out <= 4'b0000;
		 4'b0001: out <= 4'b0001;
		 4'b0010: out <= 4'b0010;
		 4'b0011: out <= 4'b0011;
		 4'b0100: out <= 4'b0100;
		 
		 //If greater than or equal to five
		 4'b0101: out <= 4'b1000;
		 4'b0110: out <= 4'b1001;
		 4'b0111: out <= 4'b1010;
		 4'b1000: out <= 4'b1011;
		 4'b1001: out <= 4'b1100;
		 4'b1010: out <= 4'b1101;
		 4'b1011: out <= 4'b1110;
		 4'b1100: out <= 4'b1111;
		
		 default: out <=4'b0000;
		
		endcase
		 
		 
endmodule
